LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY  WREG IS
PORT( 
ENTRA: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
SALE: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);   
LEER: IN STD_LOGIC;
CLKD,CLKC: IN STD_LOGIC
);
END WREG;

ARCHITECTURE NARQ OF WREG IS
BEGIN     

PROCESS (CLKD)
	BEGIN    
	IF CLKD='1'  AND CLKD'EVENT   THEN 
		IF LEER='1'  THEN  
			SALE<=ENTRA;
		END IF;
	END IF;  
	END PROCESS;                          
END NARQ;           