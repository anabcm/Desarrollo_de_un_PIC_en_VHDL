LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;   
USE IEEE.STD_LOGIC_UNSIGNED.ALL;      
USE IEEE.NUMERIC_BIT.ALL;
ENTITY RAM IS
PORT (
CLKB,CLKC,CLKD: in STD_LOGIC;
DIRECCION: in STD_LOGIC_VECTOR(8 DOWNTO 0);
BUSD: INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);   
LEER: IN STD_LOGIC;
ESCRIBIR: IN STD_LOGIC;
E_RAM:IN STD_LOGIC);
END RAM;  

ARCHITECTURE NARQ OF RAM IS
TYPE MEMORIA IS ARRAY (0 TO 511) OF STD_LOGIC_VECTOR(7 DOWNTO 0); 
SIGNAL RAM:MEMORIA;
BEGIN
PROCESS(CLKB,CLKD,CLKC)
BEGIN   
  			
 	IF(CLKB'EVENT AND CLKB='1') THEN 
			IF(ESCRIBIR='1' AND E_RAM='1') THEN
                      BUSD<=RAM(CONV_INTEGER(DIRECCION));
			ELSE
                      BUSD<="ZZZZZZZZ"; 
			END IF ;       
	ELSE

		IF(CLKD='1' AND CLKD'EVENT) THEN   
		  		IF(LEER='0' AND E_RAM='1') THEN
							  RAM(CONV_INTEGER(DIRECCION))<=BUSD;--GUARDA EL DATO     --SACA EL DATO
				END IF ;
		
      	ELSE 
			IF(CLKC='1' AND CLKC'EVENT ) THEN   
				BUSD<="ZZZZZZZZ";
			END IF;
             	 --IF(CLKB='0' AND CLKB'EVENT) THEN  BUSD<="ZZZZZZZZ"; END IF;
             	 
	 	END IF;
	END IF;	 	  

END PROCESS;
END NARQ;