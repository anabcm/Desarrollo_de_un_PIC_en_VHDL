--INTRUCTION REG
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY INS_REG IS  
PORT (     
PROGRAM_BUS:IN STD_LOGIC_VECTOR(13 DOWNTO 0);
DIRECT_ADDR:OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
DECO_BUS: OUT STD_LOGIC_VECTOR(13 DOWNTO 0); 
BIT_OPERA: OUT STD_LOGIC_VECTOR(2 DOWNTO 0); 
DIR_PC: OUT STD_LOGIC_VECTOR(10 DOWNTO 0);
CONS:OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
FLUSH: IN STD_LOGIC
);
END INS_REG;

ARCHITECTURE NARQ OF INS_REG IS
BEGIN
PROCESS (PROGRAM_BUS,FLUSH)     
	BEGIN                 
	IF(PROGRAM_BUS'EVENT) THEN
	DIRECT_ADDR<=PROGRAM_BUS(6 DOWNTO 0);
	DECO_BUS<=PROGRAM_BUS;
	BIT_OPERA<=PROGRAM_BUS(11 DOWNTO 9);
	CONS<=PROGRAM_BUS(7 DOWNTO 0);		
	ELSE
		IF(FLUSH'EVENT) THEN
			DECO_BUS<="00000000000000";  --HACE NOP EN CASO DE SER CALL O RETURN...
			
	     END IF;
  END IF;
  END PROCESS;
END NARQ;

