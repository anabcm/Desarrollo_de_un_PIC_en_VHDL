LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY DECO IS  
PORT (
   CLKA: IN STD_LOGIC;       
    BUS_ENTRA:IN STD_LOGIC_VECTOR(13 DOWNTO 0 );
    SALIDA: OUT STD_LOGIC_VECTOR(4 DOWNTO 0);   
    SD:OUT STD_LOGIC; --DICE SI HAY DIRECCIONAMIENTO INMEDIATO  
    PC,GOT:OUT STD_LOGIC;
    LEER: OUT STD_LOGIC;
    ESCRIBIR: OUT STD_LOGIC
);
END DECO;              

ARCHITECTURE NARQ OF DECO IS
BEGIN
PROCESS (CLKA)
VARIABLE CTRL: STD_LOGIC_VECTOR( 1 DOWNTO 0);  --DECODIFICADOR COMPLETO
VARIABLE FROP: STD_LOGIC_VECTOR( 1 DOWNTO 0);   --FILE REGISTER OPERATION
VARIABLE BOFR: STD_LOGIC_VECTOR( 3 DOWNTO 0);   --BYTE ORIENTED FILE REGISTER
VARIABLE LACO: STD_LOGIC_VECTOR( 2 DOWNTO 0);   --BYTE ORIENTED FILE REGISTER  
VARIABLE WR: STD_LOGIC_VECTOR( 1 DOWNTO 0);  --PARA REGISTRO DE TRABAJO         
BEGIN  
CTRL(1 DOWNTO 0):=BUS_ENTRA(13 DOWNTO 12);  
FROP(1 DOWNTO 0):=BUS_ENTRA(11 DOWNTO 10);  
BOFR(3 DOWNTO 0):=BUS_ENTRA(11 DOWNTO 8); 
LACO(2 DOWNTO 0):=BUS_ENTRA(11 DOWNTO 9);
WR(1 DOWNTO 0):=BUS_ENTRA(11 DOWNTO 10);   
PC<='U';
GOT<='0';
IF (CLKA='1') THEN               
      SD<='0';  --NADIE ESCRIBE EN EL BUS-NI LEE DEL BUS
	CASE CTRL IS
	WHEN "00" =>  	 --MANEJA UN SALIDA DE F, HABILITA EL MUX MUTANTE Y LE DICE SI PONERSE EN ALTA IMPEDANCIA O NO   
		    --CASOS DE STACK        
		    CASE BUS_ENTRA(11 DOWNTO 0) IS
			    WHEN "000000001001" =>PC<='0';--HABILITA HACE POP DE LA PILA    RETFIE
			    WHEN "000000001000" => PC<='0';-- SE HACE POP DE LA PILA RETURN
		    END CASE; 
			CASE BOFR IS
		    WHEN "0000" =>     
		    		    CASE BUS_ENTRA(7) IS
			    		WHEN '0'=>SALIDA<="00001";--ESCRIBIR<='0';LEER<='0';   
			    		WHEN '1'=>SALIDA<="00010";ESCRIBIR<='1'; IF(BUS_ENTRA(7)='1')     THEN LEER<='0';  ELSE LEER<='1';  END IF;--MOVWF
		    		END CASE;
		    		SD<='0';
		    WHEN "0001" =>
		            CASE BUS_ENTRA(7) IS
			    		WHEN '1'=>SALIDA<="00011";ESCRIBIR<='1';LEER<='0';SD<='0';   --CLRF
			    		WHEN '0'=>SALIDA<="00100";ESCRIBIR<='0';LEER<='1';   --CLRW   --101 --LE TOCA AL WREG	    		
			    	END CASE;
            WHEN "0010" =>SALIDA<="00101";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1') THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--SUBWF
            WHEN "0011" =>SALIDA<="00110";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1') THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--DECF
		    WHEN "0100" =>SALIDA<="00111";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1') THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--IORWF    
		    WHEN "0101" =>SALIDA<="01000";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1') THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--ANDWF  
		    WHEN "0110" =>SALIDA<="01001";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1') THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--XORWF  
		    WHEN "0111" =>SALIDA<="01010";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1') THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--ADDWF		     
		    WHEN "1000" =>SALIDA<="01011";ESCRIBIR<='1'; IF(BUS_ENTRA(7)='1')THEN LEER<='0';  ELSE LEER<='1';  END IF; SD<='0';--MOVF  		    
		    WHEN "1001" =>SALIDA<="01100";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1') THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--COMF
		    WHEN "1010" =>SALIDA<="01101";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1') THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--INCF
		    WHEN "1011" =>SALIDA<="01110";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1')THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--DECFSZ
            WHEN "1100" =>SALIDA<="01111";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1')THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--RRF
            WHEN "1101" =>SALIDA<="10000";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1')THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--RLF  
            WHEN "1110" =>SALIDA<="10001";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1')THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--SWAPF
            WHEN "1111" =>SALIDA<="10010";ESCRIBIR<='1';IF(BUS_ENTRA(7)='1')THEN LEER<='0';  ELSE LEER<='1';  END IF;SD<='0';--INCFSZ

		END CASE;
	       
	WHEN "01" => --HABILITA EL MUX 	
	      CASE FROP IS
		      WHEN "00"=>SALIDA<="10011";LEER<='1';ESCRIBIR<='1';SD<='0';--BCF     
		      WHEN "01"=>SALIDA<="10100";LEER<='1';ESCRIBIR<='1';SD<='0';--BSF  
		      WHEN "10"=>SALIDA<="10101";LEER<='1';ESCRIBIR<='1';SD<='0';--BTFSC 
		      WHEN "11"=>SALIDA<="10110";LEER<='1';ESCRIBIR<='1';SD<='0';--BTFSS   
	      END CASE;	       	
	WHEN "10" =>  
		CASE BUS_ENTRA(11) IS
		      WHEN '0'=>PC<='1';ESCRIBIR<='0';LEER<='0';--CALL  --     
		      WHEN '1'=>GOT<='1'; ESCRIBIR<='0';LEER<='0';--GOTO         	
		 END CASE;	  
	             SD<='1';

	WHEN "11" =>    SD<='1';--LE TOCA AL WREG
                     
		IF WR= "00" THEN SALIDA<="11110";LEER<='1'; ESCRIBIR<='0'; --MOVLW      si
		END IF;
	    CASE LACO IS
	      WHEN "111"=>SALIDA<="11001";LEER<='1'; ESCRIBIR<='0';--ADDLW si   
	      WHEN "110"=>SALIDA<="11010";LEER<='1'; ESCRIBIR<='0';--SUBLW  
	      WHEN "101"=>SALIDA<="11011";LEER<='1'; ESCRIBIR<='0';--XORLW     si
	      WHEN "100"=> 
		      CASE BUS_ENTRA(8) is
			      WHEN '0'=>SALIDA<="11100";LEER<='1'; ESCRIBIR<='0';--IORLW  
			      WHEN '1'=>SALIDA<="11101";LEER<='1'; ESCRIBIR<='0';--ANDLW
		      END CASE;	 
	      END CASE;
	          
	WHEN OTHERS => SALIDA<="00000";  
    END CASE; 
    
END IF;
END PROCESS;
END NARQ;

