LIBRARY ieee;
USE IEEE.STD_LOGIC_1164.ALL; 
USE IEEE.STD_LOGIC_UNSIGNED.ALL;    
ENTITY EPROM  is
GENERIC (
BITS: INTEGER:=8;
WORDS: INTEGER:=38
);

PORT ( 
CLKD:IN STD_LOGIC;
addr: IN STD_LOGIC_VECTOR(12 DOWNTO 0);
salida: OUT STD_LOGIC_VECTOR(13 DOWNTO 0)
);
END EPROM;

ARCHITECTURE NARS OF EPROM IS 

TYPE VECTOR_ARRAY IS ARRAY (0 TO WORDS-1) OF STD_LOGIC_VECTOR(13 DOWNTO 0);
CONSTANT memory :vector_array:=(
"00000000000000",  --0
"11000011110000",
"11111000000001",
"11000000000001",
"11100111111111",
"11100011111110", --5
"11110011111111",
"11101010101010",
"11000011110000",
"00000010100000",
"11000000000001",  --A
"00000010100001",
"11000000000010",
"00000010100010", 
"00000010100000",
"00100010100010", --F
"00011110100000",
"00100010100000",
"00010110100001",
"00000110100010",
"00000100000011",
"00100110100000",--15
"00001110100001",
"00101110100000",
"00101010100010",
"00000010100000",
"00000000000000",
"00110110100001",
"00110010100010",
"00001010100000",
"00111010100001",
"00011010100010",
"01000000100000",
"01010000100001",
"01100000100010",
"00000000000000",
"01110000100000",
"00000000000000");
BEGIN 
PROCESS (addr,CLKD)
BEGIN 
IF(CLKD ='1' AND CLKD'EVENT)  THEN
	salida<=memory(CONV_INTEGER(addr));
END IF;
END PROCESS;
end NARS;